package opcodes is
    type opcode_t is (
        OAdd,
        OSub,
        OMulH,
        OMulL,
        OShiftLeft,
        OShiftRight,
        ORotateLeft,
        ORotateRigth,
        ONot,
        OAnd,
        OOr,
        OXor,
        ODiv,
        OMod
    );
end package opcodes;

package body opcodes is

end package body opcodes;
